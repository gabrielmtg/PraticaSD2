--implementar, acho que podemos fazer isso já no somador