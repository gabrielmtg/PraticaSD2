--tem que colocar em um .do
--force /clk 0 0 ns, 1 5 ns -repeat 10 ns
--force /reset 1 0 ns, 0 10 ns
--force /enable 0 0 ns, 1 10 ns
--force /sample_ori 00000000000000000000000000000000 0 ns, 11111111111111111111111111111111 540 ns, 11111111000000001111111100000000 810 ns, 11111111000000000101010110101010 1050 ns
--force /sample_can 11111111111111111111111111111111 0 ns, 11111111111111111111111111111111 540 ns, 11111111000000001111111100000000 810 ns,  10101010010101010000000000001111 1050 ns
